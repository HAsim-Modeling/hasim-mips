import hasim_isa::*;

Addr pcStart = 32'h00001000;

typedef 4 FetchWidth;
typedef 4 CommitWidth;
typedef 32 ROBCount;
typedef 16 IntQCount;
typedef 16 MemQCount;
typedef 32 FreeListCount;
typedef 4 BranchCount;
typedef 5 NumFuncUnits;
typedef 64 PRNum;
