
import hasim_common::*;

module [HASIM_MODULE] mkMemory
    //interface:
                (Empty);

endmodule
