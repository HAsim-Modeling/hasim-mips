
import hasim_common::*;

module [HASim_Module] mkMemory
    //interface:
                (Empty);

endmodule
