import hasim_common::*;
import hasim_isa::*;

import Vector::*;

import hasim_cpu_types::*;
import hasim_cpu_parameters::*;

typedef enum {Fetch, FetchDone} FetchState deriving (Bits, Eq);

module [HASim_Module] mkPipe_Fetch();
    Connection_Send#(Bit#(8))              fpTokReq <- mkConnection_Send("fp_tok_req");
    Connection_Receive#(Token)            fpTokResp <- mkConnection_Receive("fp_tok_resp");
    Connection_Send#(Tuple2#(Token, Addr)) fpFetReq <- mkConnection_Send("fp_fet_req");

    Port_Receive#(FetchCount)        fetchCountPort <- mkPort_Receive("fetchCount", 1);
    Port_Receive#(Addr)           predictedAddrPort <- mkPort_Receive("predictedAddr", 1);
    Port_Receive#(Addr)          mispredictAddrPort <- mkPort_Receive("mispredictAddr", 1);

    Port_Send#(Addr)                   instAddrPort <- mkPort_Send("instAddr");

    Reg#(FetchState)                     fetchState <- mkReg(FetchDone);
    Reg#(Addr)                                   pc <- mkReg(pcStart);
    Reg#(FetchCount)                     totalCount <- mkReg(?);
    Reg#(FetchCount)                       fetchPos <- mkReg(?);

    Reg#(Bool)                     fillFetchInvalid <- mkReg(False);

    Reg#(ClockCounter)                     clockReg <- mkReg(0);
    Reg#(ClockCounter)                     modelReg <- mkReg(0);

    Reg#(TIMEP_Epoch)                         epoch <- mkReg(0);

    rule clockCount(True);
        clockReg <= clockReg + 1;
    endrule

    rule synchronize(fetchState == FetchDone);
        modelReg <= modelReg + 1;
        Maybe#(Addr)    predictedAddr <- predictedAddrPort.receive();
        Maybe#(Addr)   mispredictAddr <- mispredictAddrPort.receive();
        Maybe#(FetchCount) fetchCount <- fetchCountPort.receive();

        if(isValid(mispredictAddr))
        begin
            pc    <= validValue(mispredictAddr);
            epoch <= epoch + 1;
        end
        else if(isValid(predictedAddr))
        begin
            pc <= validValue(predictedAddr);
        end
        else
        begin
            pc <= pc;
        end

        FetchCount newCount = fromMaybe(fromInteger(valueOf(FetchWidth)), fetchCount);
        totalCount   <= newCount;
        fetchPos     <= 0;

        fetchState <= Fetch;

        if(newCount == 0)
        begin
            fillFetchInvalid <= True;
        end
        else
        begin
            $display("0 1 %0d %0d", clockReg, modelReg);
            fpTokReq.send(17);
            fillFetchInvalid <= False;
        end
    endrule

    rule fetch(fetchState == Fetch);
        fetchPos <= fetchPos + 1;
        if(fetchPos == fromInteger(valueOf(TSub#(FetchWidth,1))))
            fetchState <= FetchDone;
        if(!fillFetchInvalid)
        begin
            Token token <- fpTokResp.receive();
            token.timep_info = TIMEP_TokInfo{epoch: epoch,
                                             scratchpad: 0};

            fpFetReq.send(tuple2(token, pc));
            instAddrPort.send(tagged Valid pc);

            pc        <= pc + 4;
            if(fetchPos + 1 != totalCount)
                fpTokReq.send(17);
            else
                fillFetchInvalid <= True;
        end
        else
        begin
            instAddrPort.send(tagged Invalid);
        end
    endrule
endmodule
