import hasim_isa::*;

typedef 4 FetchWidth;
Addr pcStart = 32'h00001000;

typedef 32 ROBCount;
typedef 4 CommitWidth;
typedef 16 IntQCount;
typedef 16 AddrQCount;
typedef 32 FreeListCount;
typedef 4 BranchCount;
typedef 5 NumFuncUnits;
typedef 64 PRNum;
