
import hasim_base::*;
import hasim_fpgalib::*;
import hasim_common::*;

module [HASim_Module] mkMemory
    //interface:
                (Empty);

endmodule
